module BOC_PRN_GEN(rx_clk,rx_rst,
					tx_loc_boc,tx_loc_prn);

parameter ACC_WIDTH = 32;
input rx_clk,rx_rst;

output tx_loc_boc,tx_loc_prn;

